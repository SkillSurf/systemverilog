module adder32 (Ci,
    Co,
    A,
    B,
    S);
 input Ci;
 output Co;
 input [31:0] A;
 input [31:0] B;
 output [31:0] S;

 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;

 sg13g2_nand2_1 _212_ (.Y(_211_),
    .A(net57),
    .B(net25));
 sg13g2_inv_1 _213_ (.Y(_000_),
    .A(net24));
 sg13g2_nand2_2 _214_ (.Y(_001_),
    .A(net52),
    .B(net20));
 sg13g2_or2_1 _215_ (.X(_002_),
    .B(net32),
    .A(net64));
 sg13g2_inv_1 _216_ (.Y(_003_),
    .A(net63));
 sg13g2_inv_1 _217_ (.Y(_004_),
    .A(net31));
 sg13g2_nor2_1 _218_ (.A(_003_),
    .B(_004_),
    .Y(_005_));
 sg13g2_and2_1 _219_ (.A(net64),
    .B(net32),
    .X(_006_));
 sg13g2_a221oi_1 _220_ (.B2(_005_),
    .C1(_006_),
    .B1(_002_),
    .A1(net34),
    .Y(_007_),
    .A2(net2));
 sg13g2_or2_1 _221_ (.X(_008_),
    .B(net3),
    .A(net35));
 sg13g2_o21ai_1 _222_ (.B1(_008_),
    .Y(_009_),
    .A1(net34),
    .A2(net2));
 sg13g2_nand2_1 _223_ (.Y(_010_),
    .A(net35),
    .B(net3));
 sg13g2_o21ai_1 _224_ (.B1(_010_),
    .Y(_011_),
    .A1(_007_),
    .A2(_009_));
 sg13g2_xnor2_1 _225_ (.Y(_012_),
    .A(net41),
    .B(net9));
 sg13g2_xor2_1 _226_ (.B(net8),
    .A(net40),
    .X(_013_));
 sg13g2_nand2b_1 _227_ (.Y(_014_),
    .B(_013_),
    .A_N(_012_));
 sg13g2_xor2_1 _228_ (.B(net4),
    .A(net36),
    .X(_015_));
 sg13g2_xor2_1 _229_ (.B(net7),
    .A(net39),
    .X(_016_));
 sg13g2_xor2_1 _230_ (.B(net5),
    .A(net37),
    .X(_017_));
 sg13g2_xor2_1 _231_ (.B(net6),
    .A(net38),
    .X(_018_));
 sg13g2_nand4_1 _232_ (.B(_016_),
    .C(_017_),
    .A(_015_),
    .Y(_019_),
    .D(_018_));
 sg13g2_nor2_1 _233_ (.A(_014_),
    .B(_019_),
    .Y(_020_));
 sg13g2_xor2_1 _234_ (.B(net32),
    .A(net64),
    .X(_021_));
 sg13g2_xor2_1 _235_ (.B(net31),
    .A(net63),
    .X(_022_));
 sg13g2_nand2_1 _236_ (.Y(_023_),
    .A(_021_),
    .B(_022_));
 sg13g2_xor2_1 _237_ (.B(net3),
    .A(net35),
    .X(_024_));
 sg13g2_inv_1 _238_ (.Y(_025_),
    .A(_024_));
 sg13g2_xnor2_1 _239_ (.Y(_026_),
    .A(net34),
    .B(net2));
 sg13g2_or2_1 _240_ (.X(_027_),
    .B(_026_),
    .A(_025_));
 sg13g2_nor4_1 _241_ (.A(_023_),
    .B(_027_),
    .C(_014_),
    .D(_019_),
    .Y(_028_));
 sg13g2_or2_1 _242_ (.X(_029_),
    .B(net65),
    .A(net1));
 sg13g2_a21o_1 _243_ (.A2(net65),
    .A1(net1),
    .B1(net33),
    .X(_030_));
 sg13g2_a22oi_1 _244_ (.Y(_031_),
    .B1(_029_),
    .B2(_030_),
    .A2(net12),
    .A1(net44));
 sg13g2_nor2_1 _245_ (.A(net44),
    .B(net12),
    .Y(_032_));
 sg13g2_xor2_1 _246_ (.B(net26),
    .A(net58),
    .X(_033_));
 sg13g2_xor2_1 _247_ (.B(net23),
    .A(net55),
    .X(_034_));
 sg13g2_nand3b_1 _248_ (.B(_033_),
    .C(_034_),
    .Y(_035_),
    .A_N(_032_));
 sg13g2_nor2_1 _249_ (.A(net58),
    .B(net26),
    .Y(_036_));
 sg13g2_a22oi_1 _250_ (.Y(_037_),
    .B1(net58),
    .B2(net26),
    .A2(net23),
    .A1(net55));
 sg13g2_or2_1 _251_ (.X(_038_),
    .B(_037_),
    .A(_036_));
 sg13g2_o21ai_1 _252_ (.B1(_038_),
    .Y(_039_),
    .A1(_031_),
    .A2(_035_));
 sg13g2_xor2_1 _253_ (.B(net28),
    .A(net60),
    .X(_040_));
 sg13g2_xor2_1 _254_ (.B(net27),
    .A(net59),
    .X(_041_));
 sg13g2_nand2_1 _255_ (.Y(_042_),
    .A(_040_),
    .B(_041_));
 sg13g2_xor2_1 _256_ (.B(net30),
    .A(net62),
    .X(_043_));
 sg13g2_xor2_1 _257_ (.B(net29),
    .A(net61),
    .X(_044_));
 sg13g2_nand2_1 _258_ (.Y(_045_),
    .A(_043_),
    .B(_044_));
 sg13g2_nor2_1 _259_ (.A(_042_),
    .B(_045_),
    .Y(_046_));
 sg13g2_or2_1 _260_ (.X(_047_),
    .B(net28),
    .A(net60));
 sg13g2_and2_1 _261_ (.A(net59),
    .B(net27),
    .X(_048_));
 sg13g2_and2_1 _262_ (.A(net60),
    .B(net28),
    .X(_049_));
 sg13g2_a221oi_1 _263_ (.B2(_048_),
    .C1(_049_),
    .B1(_047_),
    .A1(net61),
    .Y(_050_),
    .A2(net29));
 sg13g2_or2_1 _264_ (.X(_051_),
    .B(net30),
    .A(net62));
 sg13g2_o21ai_1 _265_ (.B1(_051_),
    .Y(_052_),
    .A1(net61),
    .A2(net29));
 sg13g2_nand2_1 _266_ (.Y(_053_),
    .A(net62),
    .B(net30));
 sg13g2_o21ai_1 _267_ (.B1(_053_),
    .Y(_054_),
    .A1(_050_),
    .A2(_052_));
 sg13g2_a21o_1 _268_ (.A2(_046_),
    .A1(_039_),
    .B1(_054_),
    .X(_055_));
 sg13g2_a22oi_1 _269_ (.Y(_056_),
    .B1(_028_),
    .B2(_055_),
    .A2(_020_),
    .A1(_011_));
 sg13g2_or2_1 _270_ (.X(_057_),
    .B(net9),
    .A(net41));
 sg13g2_and3_1 _271_ (.X(_058_),
    .A(net40),
    .B(net8),
    .C(_057_));
 sg13g2_a21oi_1 _272_ (.A1(net41),
    .A2(net9),
    .Y(_059_),
    .B1(_058_));
 sg13g2_inv_1 _273_ (.Y(_060_),
    .A(_059_));
 sg13g2_or2_1 _274_ (.X(_061_),
    .B(net6),
    .A(net38));
 sg13g2_nand2_1 _275_ (.Y(_062_),
    .A(net36),
    .B(net4));
 sg13g2_nor2_1 _276_ (.A(net37),
    .B(net5),
    .Y(_063_));
 sg13g2_a22oi_1 _277_ (.Y(_064_),
    .B1(net38),
    .B2(net6),
    .A2(net5),
    .A1(net37));
 sg13g2_o21ai_1 _278_ (.B1(_064_),
    .Y(_065_),
    .A1(_062_),
    .A2(_063_));
 sg13g2_a22oi_1 _279_ (.Y(_066_),
    .B1(_061_),
    .B2(_065_),
    .A2(net7),
    .A1(net39));
 sg13g2_nor2_1 _280_ (.A(net39),
    .B(net7),
    .Y(_067_));
 sg13g2_o21ai_1 _281_ (.B1(_057_),
    .Y(_068_),
    .A1(net40),
    .A2(net8));
 sg13g2_nor3_1 _282_ (.A(_066_),
    .B(_067_),
    .C(_068_),
    .Y(_069_));
 sg13g2_nor2_1 _283_ (.A(net43),
    .B(net11),
    .Y(_070_));
 sg13g2_nand2_1 _284_ (.Y(_071_),
    .A(net42),
    .B(net10));
 sg13g2_nand2_1 _285_ (.Y(_072_),
    .A(net43),
    .B(net11));
 sg13g2_o21ai_1 _286_ (.B1(_072_),
    .Y(_073_),
    .A1(_070_),
    .A2(_071_));
 sg13g2_nor2_1 _287_ (.A(net46),
    .B(net14),
    .Y(_074_));
 sg13g2_nand2_1 _288_ (.Y(_075_),
    .A(net45),
    .B(net13));
 sg13g2_nand2_1 _289_ (.Y(_076_),
    .A(net46),
    .B(net14));
 sg13g2_o21ai_1 _290_ (.B1(_076_),
    .Y(_077_),
    .A1(_074_),
    .A2(_075_));
 sg13g2_nor4_1 _291_ (.A(_060_),
    .B(_069_),
    .C(_073_),
    .D(_077_),
    .Y(_078_));
 sg13g2_xnor2_1 _292_ (.Y(_079_),
    .A(net43),
    .B(net11));
 sg13g2_xnor2_1 _293_ (.Y(_080_),
    .A(net42),
    .B(net10));
 sg13g2_nor2_1 _294_ (.A(_079_),
    .B(_080_),
    .Y(_081_));
 sg13g2_or2_1 _295_ (.X(_082_),
    .B(_073_),
    .A(_081_));
 sg13g2_nor2_1 _296_ (.A(net45),
    .B(net13),
    .Y(_083_));
 sg13g2_a21oi_1 _297_ (.A1(_083_),
    .A2(_076_),
    .Y(_084_),
    .B1(_074_));
 sg13g2_o21ai_1 _298_ (.B1(_084_),
    .Y(_085_),
    .A1(_077_),
    .A2(_082_));
 sg13g2_a21oi_2 _299_ (.B1(_085_),
    .Y(_086_),
    .A2(_078_),
    .A1(_056_));
 sg13g2_nor2_1 _300_ (.A(net50),
    .B(net18),
    .Y(_087_));
 sg13g2_a22oi_1 _301_ (.Y(_088_),
    .B1(net50),
    .B2(net18),
    .A2(net17),
    .A1(net49));
 sg13g2_nor2_1 _302_ (.A(_087_),
    .B(_088_),
    .Y(_089_));
 sg13g2_nor2_1 _303_ (.A(net19),
    .B(_089_),
    .Y(_090_));
 sg13g2_nand2_1 _304_ (.Y(_091_),
    .A(net47),
    .B(net15));
 sg13g2_or2_1 _305_ (.X(_092_),
    .B(net16),
    .A(net48));
 sg13g2_nor2b_1 _306_ (.A(_091_),
    .B_N(_092_),
    .Y(_093_));
 sg13g2_a21oi_2 _307_ (.B1(_093_),
    .Y(_094_),
    .A2(net16),
    .A1(net48));
 sg13g2_nand2_1 _308_ (.Y(_095_),
    .A(_090_),
    .B(_094_));
 sg13g2_xor2_1 _309_ (.B(net16),
    .A(net48),
    .X(_096_));
 sg13g2_xor2_1 _310_ (.B(net15),
    .A(net47),
    .X(_097_));
 sg13g2_nand2_1 _311_ (.Y(_098_),
    .A(_096_),
    .B(_097_));
 sg13g2_xor2_1 _312_ (.B(net18),
    .A(net50),
    .X(_099_));
 sg13g2_xor2_1 _313_ (.B(net17),
    .A(net49),
    .X(_100_));
 sg13g2_nand2_1 _314_ (.Y(_101_),
    .A(_099_),
    .B(_100_));
 sg13g2_a21o_1 _315_ (.A2(_098_),
    .A1(_094_),
    .B1(_101_),
    .X(_102_));
 sg13g2_nor2_1 _316_ (.A(net52),
    .B(net20),
    .Y(_103_));
 sg13g2_a21oi_1 _317_ (.A1(_090_),
    .A2(_102_),
    .Y(_104_),
    .B1(_103_));
 sg13g2_o21ai_1 _318_ (.B1(_104_),
    .Y(_105_),
    .A1(_086_),
    .A2(_095_));
 sg13g2_nand2_1 _319_ (.Y(_106_),
    .A(net21),
    .B(net54));
 sg13g2_nand2_1 _320_ (.Y(_107_),
    .A(net53),
    .B(net54));
 sg13g2_inv_1 _321_ (.Y(_108_),
    .A(net19));
 sg13g2_nor3_1 _322_ (.A(_108_),
    .B(_101_),
    .C(_098_),
    .Y(_109_));
 sg13g2_nor2_1 _323_ (.A(_101_),
    .B(_094_),
    .Y(_110_));
 sg13g2_o21ai_1 _324_ (.B1(net19),
    .Y(_111_),
    .A1(_089_),
    .A2(_110_));
 sg13g2_nand3b_1 _325_ (.B(_001_),
    .C(_111_),
    .Y(_112_),
    .A_N(net51));
 sg13g2_a21oi_2 _326_ (.B1(_112_),
    .Y(_113_),
    .A2(_109_),
    .A1(_086_));
 sg13g2_a221oi_1 _327_ (.B2(_107_),
    .C1(_113_),
    .B1(_106_),
    .A1(_001_),
    .Y(_114_),
    .A2(_105_));
 sg13g2_nand2_1 _328_ (.Y(_115_),
    .A(net21),
    .B(net22));
 sg13g2_nand2_1 _329_ (.Y(_116_),
    .A(net53),
    .B(net22));
 sg13g2_a221oi_1 _330_ (.B2(_116_),
    .C1(_113_),
    .B1(_115_),
    .A1(_001_),
    .Y(_117_),
    .A2(_105_));
 sg13g2_or2_1 _331_ (.X(_118_),
    .B(net22),
    .A(net54));
 sg13g2_nand3_1 _332_ (.B(net21),
    .C(_118_),
    .A(net53),
    .Y(_119_));
 sg13g2_nand2_1 _333_ (.Y(_120_),
    .A(net54),
    .B(net22));
 sg13g2_nand2_1 _334_ (.Y(_121_),
    .A(_119_),
    .B(_120_));
 sg13g2_nor3_1 _335_ (.A(_114_),
    .B(_117_),
    .C(_121_),
    .Y(_122_));
 sg13g2_nand3_1 _336_ (.B(net24),
    .C(_118_),
    .A(net21),
    .Y(_123_));
 sg13g2_nand3_1 _337_ (.B(net24),
    .C(_118_),
    .A(net53),
    .Y(_124_));
 sg13g2_a221oi_1 _338_ (.B2(_124_),
    .C1(_113_),
    .B1(_123_),
    .A1(_001_),
    .Y(_125_),
    .A2(_105_));
 sg13g2_a21oi_1 _339_ (.A1(_119_),
    .A2(_120_),
    .Y(_126_),
    .B1(_000_));
 sg13g2_nor3_1 _340_ (.A(net56),
    .B(_125_),
    .C(_126_),
    .Y(_127_));
 sg13g2_a21o_1 _341_ (.A2(_122_),
    .A1(_000_),
    .B1(_127_),
    .X(_128_));
 sg13g2_nor2_1 _342_ (.A(net57),
    .B(net25),
    .Y(_129_));
 sg13g2_a21oi_1 _343_ (.A1(_211_),
    .A2(_128_),
    .Y(net66),
    .B1(_129_));
 sg13g2_xnor2_1 _344_ (.Y(_130_),
    .A(net1),
    .B(net65));
 sg13g2_xnor2_1 _345_ (.Y(net67),
    .A(net33),
    .B(_130_));
 sg13g2_nand3_1 _346_ (.B(net29),
    .C(_051_),
    .A(net61),
    .Y(_131_));
 sg13g2_a22oi_1 _347_ (.Y(_132_),
    .B1(_053_),
    .B2(_131_),
    .A2(_004_),
    .A1(_003_));
 sg13g2_or2_1 _348_ (.X(_133_),
    .B(_132_),
    .A(_005_));
 sg13g2_a21oi_1 _349_ (.A1(net32),
    .A2(_133_),
    .Y(_134_),
    .B1(net64));
 sg13g2_nor2_1 _350_ (.A(net32),
    .B(_133_),
    .Y(_135_));
 sg13g2_inv_1 _351_ (.Y(_136_),
    .A(_042_));
 sg13g2_a221oi_1 _352_ (.B2(_136_),
    .C1(_049_),
    .B1(_039_),
    .A1(_047_),
    .Y(_137_),
    .A2(_048_));
 sg13g2_or3_1 _353_ (.A(_045_),
    .B(_023_),
    .C(_137_),
    .X(_138_));
 sg13g2_o21ai_1 _354_ (.B1(_138_),
    .Y(_139_),
    .A1(_134_),
    .A2(_135_));
 sg13g2_xnor2_1 _355_ (.Y(net68),
    .A(_026_),
    .B(_139_));
 sg13g2_a21o_1 _356_ (.A2(_139_),
    .A1(net2),
    .B1(net34),
    .X(_140_));
 sg13g2_o21ai_1 _357_ (.B1(_140_),
    .Y(_141_),
    .A1(net2),
    .A2(_139_));
 sg13g2_xnor2_1 _358_ (.Y(net69),
    .A(_024_),
    .B(_141_));
 sg13g2_nor2_1 _359_ (.A(_023_),
    .B(_027_),
    .Y(_142_));
 sg13g2_a21oi_2 _360_ (.B1(_011_),
    .Y(_143_),
    .A2(_142_),
    .A1(_055_));
 sg13g2_xnor2_1 _361_ (.Y(net70),
    .A(_143_),
    .B(_015_));
 sg13g2_nor2_1 _362_ (.A(net36),
    .B(net4),
    .Y(_144_));
 sg13g2_a21oi_1 _363_ (.A1(_143_),
    .A2(_062_),
    .Y(_145_),
    .B1(_144_));
 sg13g2_xor2_1 _364_ (.B(_145_),
    .A(_017_),
    .X(net71));
 sg13g2_a21o_1 _365_ (.A2(_145_),
    .A1(net5),
    .B1(net37),
    .X(_146_));
 sg13g2_o21ai_1 _366_ (.B1(_146_),
    .Y(_147_),
    .A1(net5),
    .A2(_145_));
 sg13g2_xnor2_1 _367_ (.Y(net72),
    .A(_018_),
    .B(_147_));
 sg13g2_nor2b_1 _368_ (.A(_147_),
    .B_N(_061_),
    .Y(_148_));
 sg13g2_a21oi_1 _369_ (.A1(net38),
    .A2(net6),
    .Y(_149_),
    .B1(_148_));
 sg13g2_xnor2_1 _370_ (.Y(net73),
    .A(_016_),
    .B(_149_));
 sg13g2_nor2_1 _371_ (.A(_143_),
    .B(_019_),
    .Y(_150_));
 sg13g2_nor2_1 _372_ (.A(_066_),
    .B(_067_),
    .Y(_151_));
 sg13g2_nor2_1 _373_ (.A(_150_),
    .B(_151_),
    .Y(_152_));
 sg13g2_xnor2_1 _374_ (.Y(net74),
    .A(_013_),
    .B(_152_));
 sg13g2_nor2b_1 _375_ (.A(_152_),
    .B_N(net8),
    .Y(_153_));
 sg13g2_nand2b_1 _376_ (.Y(_154_),
    .B(_152_),
    .A_N(net8));
 sg13g2_o21ai_1 _377_ (.B1(_154_),
    .Y(_155_),
    .A1(net40),
    .A2(_153_));
 sg13g2_xor2_1 _378_ (.B(_155_),
    .A(_012_),
    .X(net75));
 sg13g2_nor2_1 _379_ (.A(_060_),
    .B(_069_),
    .Y(_156_));
 sg13g2_nand2_2 _380_ (.Y(_157_),
    .A(_056_),
    .B(_156_));
 sg13g2_xnor2_1 _381_ (.Y(net76),
    .A(_157_),
    .B(_080_));
 sg13g2_o21ai_1 _382_ (.B1(_157_),
    .Y(_158_),
    .A1(net42),
    .A2(net10));
 sg13g2_nand2_1 _383_ (.Y(_159_),
    .A(_071_),
    .B(_158_));
 sg13g2_xnor2_1 _384_ (.Y(net77),
    .A(_079_),
    .B(_159_));
 sg13g2_nand2_1 _385_ (.Y(_160_),
    .A(_029_),
    .B(_030_));
 sg13g2_xor2_1 _386_ (.B(net12),
    .A(net44),
    .X(_161_));
 sg13g2_xnor2_1 _387_ (.Y(net78),
    .A(_160_),
    .B(_161_));
 sg13g2_a21oi_1 _388_ (.A1(_157_),
    .A2(_081_),
    .Y(_162_),
    .B1(_073_));
 sg13g2_xor2_1 _389_ (.B(net13),
    .A(net45),
    .X(_163_));
 sg13g2_xnor2_1 _390_ (.Y(net79),
    .A(_162_),
    .B(_163_));
 sg13g2_a221oi_1 _391_ (.B2(_081_),
    .C1(_073_),
    .B1(_157_),
    .A1(net45),
    .Y(_164_),
    .A2(net13));
 sg13g2_or2_1 _392_ (.X(_165_),
    .B(_164_),
    .A(_083_));
 sg13g2_xor2_1 _393_ (.B(net14),
    .A(net46),
    .X(_166_));
 sg13g2_xnor2_1 _394_ (.Y(net80),
    .A(_165_),
    .B(_166_));
 sg13g2_xor2_1 _395_ (.B(_086_),
    .A(_097_),
    .X(net81));
 sg13g2_nor2_1 _396_ (.A(net47),
    .B(net15),
    .Y(_167_));
 sg13g2_a21oi_1 _397_ (.A1(_091_),
    .A2(_076_),
    .Y(_168_),
    .B1(_167_));
 sg13g2_nand2_1 _398_ (.Y(_169_),
    .A(_097_),
    .B(_166_));
 sg13g2_nor2_1 _399_ (.A(_165_),
    .B(_169_),
    .Y(_170_));
 sg13g2_nor2_1 _400_ (.A(_168_),
    .B(_170_),
    .Y(_171_));
 sg13g2_xnor2_1 _401_ (.Y(net82),
    .A(_096_),
    .B(_171_));
 sg13g2_nand2b_1 _402_ (.Y(_172_),
    .B(_086_),
    .A_N(_098_));
 sg13g2_and2_1 _403_ (.A(_094_),
    .B(_172_),
    .X(_173_));
 sg13g2_xnor2_1 _404_ (.Y(net83),
    .A(_100_),
    .B(_173_));
 sg13g2_nand2b_1 _405_ (.Y(_174_),
    .B(_173_),
    .A_N(net17));
 sg13g2_nor2b_1 _406_ (.A(_173_),
    .B_N(net17),
    .Y(_175_));
 sg13g2_a21oi_1 _407_ (.A1(net49),
    .A2(_174_),
    .Y(_176_),
    .B1(_175_));
 sg13g2_xnor2_1 _408_ (.Y(net84),
    .A(_099_),
    .B(_176_));
 sg13g2_nor2_1 _409_ (.A(_101_),
    .B(_173_),
    .Y(_177_));
 sg13g2_nor2_1 _410_ (.A(_089_),
    .B(_177_),
    .Y(_178_));
 sg13g2_xor2_1 _411_ (.B(net19),
    .A(net51),
    .X(_179_));
 sg13g2_xnor2_1 _412_ (.Y(net85),
    .A(_178_),
    .B(_179_));
 sg13g2_a221oi_1 _413_ (.B2(net17),
    .C1(_168_),
    .B1(net49),
    .A1(net48),
    .Y(_180_),
    .A2(net16));
 sg13g2_o21ai_1 _414_ (.B1(_180_),
    .Y(_181_),
    .A1(_165_),
    .A2(_169_));
 sg13g2_nor2_1 _415_ (.A(net51),
    .B(net19),
    .Y(_182_));
 sg13g2_o21ai_1 _416_ (.B1(_092_),
    .Y(_183_),
    .A1(net49),
    .A2(net17));
 sg13g2_inv_1 _417_ (.Y(_184_),
    .A(_183_));
 sg13g2_a21oi_1 _418_ (.A1(net49),
    .A2(net17),
    .Y(_185_),
    .B1(_184_));
 sg13g2_nor3_1 _419_ (.A(_087_),
    .B(_182_),
    .C(_185_),
    .Y(_186_));
 sg13g2_a22oi_1 _420_ (.Y(_187_),
    .B1(net51),
    .B2(net19),
    .A2(net18),
    .A1(net50));
 sg13g2_nor2_1 _421_ (.A(_182_),
    .B(_187_),
    .Y(_188_));
 sg13g2_a21oi_1 _422_ (.A1(_181_),
    .A2(_186_),
    .Y(_189_),
    .B1(_188_));
 sg13g2_xor2_1 _423_ (.B(net20),
    .A(net52),
    .X(_190_));
 sg13g2_xnor2_1 _424_ (.Y(net86),
    .A(_189_),
    .B(_190_));
 sg13g2_a21oi_2 _425_ (.B1(_113_),
    .Y(_191_),
    .A2(_105_),
    .A1(_001_));
 sg13g2_xnor2_1 _426_ (.Y(_192_),
    .A(net53),
    .B(net21));
 sg13g2_xnor2_1 _427_ (.Y(net87),
    .A(_191_),
    .B(_192_));
 sg13g2_a21o_1 _428_ (.A2(_191_),
    .A1(net21),
    .B1(net53),
    .X(_193_));
 sg13g2_o21ai_1 _429_ (.B1(_193_),
    .Y(_194_),
    .A1(net21),
    .A2(_191_));
 sg13g2_xor2_1 _430_ (.B(net22),
    .A(net54),
    .X(_195_));
 sg13g2_xnor2_1 _431_ (.Y(net88),
    .A(_194_),
    .B(_195_));
 sg13g2_nor2_1 _432_ (.A(_031_),
    .B(_032_),
    .Y(_196_));
 sg13g2_xor2_1 _433_ (.B(_196_),
    .A(_034_),
    .X(net89));
 sg13g2_xor2_1 _434_ (.B(net24),
    .A(net56),
    .X(_197_));
 sg13g2_xnor2_1 _435_ (.Y(net90),
    .A(_122_),
    .B(_197_));
 sg13g2_xor2_1 _436_ (.B(net25),
    .A(net57),
    .X(_198_));
 sg13g2_xnor2_1 _437_ (.Y(net91),
    .A(_128_),
    .B(_198_));
 sg13g2_nor2_1 _438_ (.A(net23),
    .B(_196_),
    .Y(_199_));
 sg13g2_a21oi_1 _439_ (.A1(net23),
    .A2(_196_),
    .Y(_200_),
    .B1(net55));
 sg13g2_nor2_1 _440_ (.A(_199_),
    .B(_200_),
    .Y(_201_));
 sg13g2_xor2_1 _441_ (.B(_201_),
    .A(_033_),
    .X(net92));
 sg13g2_xor2_1 _442_ (.B(_041_),
    .A(_039_),
    .X(net93));
 sg13g2_a21oi_1 _443_ (.A1(net27),
    .A2(_039_),
    .Y(_202_),
    .B1(net59));
 sg13g2_nor2_1 _444_ (.A(net27),
    .B(_039_),
    .Y(_203_));
 sg13g2_nor2_1 _445_ (.A(_202_),
    .B(_203_),
    .Y(_204_));
 sg13g2_xor2_1 _446_ (.B(_204_),
    .A(_040_),
    .X(net94));
 sg13g2_xnor2_1 _447_ (.Y(net95),
    .A(_044_),
    .B(_137_));
 sg13g2_nand2b_1 _448_ (.Y(_205_),
    .B(_137_),
    .A_N(net29));
 sg13g2_nor2b_1 _449_ (.A(_137_),
    .B_N(net29),
    .Y(_206_));
 sg13g2_a21oi_1 _450_ (.A1(net61),
    .A2(_205_),
    .Y(_207_),
    .B1(_206_));
 sg13g2_xnor2_1 _451_ (.Y(net96),
    .A(_043_),
    .B(_207_));
 sg13g2_a21oi_1 _452_ (.A1(_039_),
    .A2(_046_),
    .Y(_208_),
    .B1(_054_));
 sg13g2_xnor2_1 _453_ (.Y(net97),
    .A(_208_),
    .B(_022_));
 sg13g2_a21oi_1 _454_ (.A1(net31),
    .A2(_055_),
    .Y(_209_),
    .B1(net63));
 sg13g2_a21oi_1 _455_ (.A1(_004_),
    .A2(_208_),
    .Y(_210_),
    .B1(_209_));
 sg13g2_xor2_1 _456_ (.B(_210_),
    .A(_021_),
    .X(net98));
 sg13g2_buf_1 input1 (.A(A[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(A[10]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(A[11]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(A[12]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(A[13]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(A[14]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(A[15]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(A[16]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(A[17]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(A[18]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(A[19]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(A[1]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(A[20]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(A[21]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(A[22]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(A[23]),
    .X(net16));
 sg13g2_buf_2 input17 (.A(A[24]),
    .X(net17));
 sg13g2_buf_1 input18 (.A(A[25]),
    .X(net18));
 sg13g2_buf_2 input19 (.A(A[26]),
    .X(net19));
 sg13g2_buf_1 input20 (.A(A[27]),
    .X(net20));
 sg13g2_buf_2 input21 (.A(A[28]),
    .X(net21));
 sg13g2_buf_1 input22 (.A(A[29]),
    .X(net22));
 sg13g2_buf_1 input23 (.A(A[2]),
    .X(net23));
 sg13g2_buf_1 input24 (.A(A[30]),
    .X(net24));
 sg13g2_buf_1 input25 (.A(A[31]),
    .X(net25));
 sg13g2_buf_1 input26 (.A(A[3]),
    .X(net26));
 sg13g2_buf_1 input27 (.A(A[4]),
    .X(net27));
 sg13g2_buf_1 input28 (.A(A[5]),
    .X(net28));
 sg13g2_buf_1 input29 (.A(A[6]),
    .X(net29));
 sg13g2_buf_1 input30 (.A(A[7]),
    .X(net30));
 sg13g2_buf_1 input31 (.A(A[8]),
    .X(net31));
 sg13g2_buf_1 input32 (.A(A[9]),
    .X(net32));
 sg13g2_buf_1 input33 (.A(B[0]),
    .X(net33));
 sg13g2_buf_1 input34 (.A(B[10]),
    .X(net34));
 sg13g2_buf_1 input35 (.A(B[11]),
    .X(net35));
 sg13g2_buf_1 input36 (.A(B[12]),
    .X(net36));
 sg13g2_buf_1 input37 (.A(B[13]),
    .X(net37));
 sg13g2_buf_1 input38 (.A(B[14]),
    .X(net38));
 sg13g2_buf_1 input39 (.A(B[15]),
    .X(net39));
 sg13g2_buf_1 input40 (.A(B[16]),
    .X(net40));
 sg13g2_buf_1 input41 (.A(B[17]),
    .X(net41));
 sg13g2_buf_1 input42 (.A(B[18]),
    .X(net42));
 sg13g2_buf_1 input43 (.A(B[19]),
    .X(net43));
 sg13g2_buf_1 input44 (.A(B[1]),
    .X(net44));
 sg13g2_buf_1 input45 (.A(B[20]),
    .X(net45));
 sg13g2_buf_1 input46 (.A(B[21]),
    .X(net46));
 sg13g2_buf_1 input47 (.A(B[22]),
    .X(net47));
 sg13g2_buf_1 input48 (.A(B[23]),
    .X(net48));
 sg13g2_buf_2 input49 (.A(B[24]),
    .X(net49));
 sg13g2_buf_1 input50 (.A(B[25]),
    .X(net50));
 sg13g2_buf_1 input51 (.A(B[26]),
    .X(net51));
 sg13g2_buf_1 input52 (.A(B[27]),
    .X(net52));
 sg13g2_buf_1 input53 (.A(B[28]),
    .X(net53));
 sg13g2_buf_1 input54 (.A(B[29]),
    .X(net54));
 sg13g2_buf_1 input55 (.A(B[2]),
    .X(net55));
 sg13g2_buf_1 input56 (.A(B[30]),
    .X(net56));
 sg13g2_buf_1 input57 (.A(B[31]),
    .X(net57));
 sg13g2_buf_1 input58 (.A(B[3]),
    .X(net58));
 sg13g2_buf_1 input59 (.A(B[4]),
    .X(net59));
 sg13g2_buf_1 input60 (.A(B[5]),
    .X(net60));
 sg13g2_buf_1 input61 (.A(B[6]),
    .X(net61));
 sg13g2_buf_1 input62 (.A(B[7]),
    .X(net62));
 sg13g2_buf_1 input63 (.A(B[8]),
    .X(net63));
 sg13g2_buf_1 input64 (.A(B[9]),
    .X(net64));
 sg13g2_buf_1 input65 (.A(Ci),
    .X(net65));
 sg13g2_buf_1 output66 (.A(net66),
    .X(Co));
 sg13g2_buf_1 output67 (.A(net67),
    .X(S[0]));
 sg13g2_buf_1 output68 (.A(net68),
    .X(S[10]));
 sg13g2_buf_1 output69 (.A(net69),
    .X(S[11]));
 sg13g2_buf_1 output70 (.A(net70),
    .X(S[12]));
 sg13g2_buf_1 output71 (.A(net71),
    .X(S[13]));
 sg13g2_buf_1 output72 (.A(net72),
    .X(S[14]));
 sg13g2_buf_1 output73 (.A(net73),
    .X(S[15]));
 sg13g2_buf_1 output74 (.A(net74),
    .X(S[16]));
 sg13g2_buf_1 output75 (.A(net75),
    .X(S[17]));
 sg13g2_buf_1 output76 (.A(net76),
    .X(S[18]));
 sg13g2_buf_1 output77 (.A(net77),
    .X(S[19]));
 sg13g2_buf_1 output78 (.A(net78),
    .X(S[1]));
 sg13g2_buf_1 output79 (.A(net79),
    .X(S[20]));
 sg13g2_buf_1 output80 (.A(net80),
    .X(S[21]));
 sg13g2_buf_1 output81 (.A(net81),
    .X(S[22]));
 sg13g2_buf_1 output82 (.A(net82),
    .X(S[23]));
 sg13g2_buf_1 output83 (.A(net83),
    .X(S[24]));
 sg13g2_buf_1 output84 (.A(net84),
    .X(S[25]));
 sg13g2_buf_1 output85 (.A(net85),
    .X(S[26]));
 sg13g2_buf_1 output86 (.A(net86),
    .X(S[27]));
 sg13g2_buf_1 output87 (.A(net87),
    .X(S[28]));
 sg13g2_buf_1 output88 (.A(net88),
    .X(S[29]));
 sg13g2_buf_1 output89 (.A(net89),
    .X(S[2]));
 sg13g2_buf_1 output90 (.A(net90),
    .X(S[30]));
 sg13g2_buf_1 output91 (.A(net91),
    .X(S[31]));
 sg13g2_buf_1 output92 (.A(net92),
    .X(S[3]));
 sg13g2_buf_1 output93 (.A(net93),
    .X(S[4]));
 sg13g2_buf_1 output94 (.A(net94),
    .X(S[5]));
 sg13g2_buf_1 output95 (.A(net95),
    .X(S[6]));
 sg13g2_buf_1 output96 (.A(net96),
    .X(S[7]));
 sg13g2_buf_1 output97 (.A(net97),
    .X(S[8]));
 sg13g2_buf_1 output98 (.A(net98),
    .X(S[9]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_4 FILLER_0_14 ();
 sg13g2_fill_2 FILLER_0_38 ();
 sg13g2_fill_1 FILLER_0_40 ();
 sg13g2_fill_2 FILLER_0_57 ();
 sg13g2_decap_4 FILLER_0_63 ();
 sg13g2_fill_2 FILLER_0_67 ();
 sg13g2_decap_4 FILLER_0_81 ();
 sg13g2_fill_2 FILLER_0_89 ();
 sg13g2_decap_8 FILLER_0_99 ();
 sg13g2_decap_8 FILLER_0_106 ();
 sg13g2_decap_8 FILLER_0_113 ();
 sg13g2_decap_8 FILLER_0_120 ();
 sg13g2_decap_8 FILLER_0_127 ();
 sg13g2_decap_8 FILLER_0_134 ();
 sg13g2_decap_8 FILLER_0_141 ();
 sg13g2_decap_8 FILLER_0_148 ();
 sg13g2_decap_8 FILLER_0_155 ();
 sg13g2_decap_4 FILLER_0_162 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_4 FILLER_1_28 ();
 sg13g2_fill_1 FILLER_1_32 ();
 sg13g2_decap_8 FILLER_1_41 ();
 sg13g2_decap_4 FILLER_1_48 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_4 FILLER_1_70 ();
 sg13g2_fill_2 FILLER_1_74 ();
 sg13g2_fill_2 FILLER_1_80 ();
 sg13g2_fill_1 FILLER_1_82 ();
 sg13g2_fill_2 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_97 ();
 sg13g2_decap_8 FILLER_1_104 ();
 sg13g2_decap_8 FILLER_1_111 ();
 sg13g2_decap_8 FILLER_1_118 ();
 sg13g2_decap_8 FILLER_1_125 ();
 sg13g2_decap_8 FILLER_1_132 ();
 sg13g2_decap_8 FILLER_1_139 ();
 sg13g2_decap_8 FILLER_1_146 ();
 sg13g2_decap_8 FILLER_1_153 ();
 sg13g2_decap_4 FILLER_1_160 ();
 sg13g2_fill_2 FILLER_1_164 ();
 sg13g2_decap_4 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_4 ();
 sg13g2_fill_2 FILLER_2_10 ();
 sg13g2_decap_4 FILLER_2_16 ();
 sg13g2_fill_2 FILLER_2_20 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_4 FILLER_2_161 ();
 sg13g2_fill_1 FILLER_2_165 ();
 sg13g2_fill_2 FILLER_3_12 ();
 sg13g2_fill_1 FILLER_3_14 ();
 sg13g2_fill_1 FILLER_3_25 ();
 sg13g2_fill_1 FILLER_3_31 ();
 sg13g2_fill_2 FILLER_3_40 ();
 sg13g2_fill_2 FILLER_3_50 ();
 sg13g2_fill_1 FILLER_3_52 ();
 sg13g2_decap_4 FILLER_3_61 ();
 sg13g2_fill_2 FILLER_3_65 ();
 sg13g2_decap_8 FILLER_3_75 ();
 sg13g2_decap_8 FILLER_3_82 ();
 sg13g2_decap_8 FILLER_3_89 ();
 sg13g2_decap_8 FILLER_3_96 ();
 sg13g2_decap_8 FILLER_3_103 ();
 sg13g2_decap_8 FILLER_3_110 ();
 sg13g2_decap_8 FILLER_3_117 ();
 sg13g2_decap_8 FILLER_3_124 ();
 sg13g2_decap_8 FILLER_3_131 ();
 sg13g2_decap_8 FILLER_3_138 ();
 sg13g2_decap_8 FILLER_3_145 ();
 sg13g2_decap_8 FILLER_3_152 ();
 sg13g2_decap_8 FILLER_3_159 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_7 ();
 sg13g2_fill_1 FILLER_4_9 ();
 sg13g2_fill_1 FILLER_4_14 ();
 sg13g2_fill_2 FILLER_4_23 ();
 sg13g2_fill_2 FILLER_4_33 ();
 sg13g2_fill_1 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_43 ();
 sg13g2_fill_2 FILLER_4_50 ();
 sg13g2_fill_2 FILLER_4_61 ();
 sg13g2_fill_1 FILLER_4_63 ();
 sg13g2_fill_2 FILLER_4_74 ();
 sg13g2_fill_1 FILLER_4_76 ();
 sg13g2_decap_8 FILLER_4_85 ();
 sg13g2_decap_8 FILLER_4_92 ();
 sg13g2_decap_8 FILLER_4_99 ();
 sg13g2_decap_8 FILLER_4_106 ();
 sg13g2_decap_8 FILLER_4_113 ();
 sg13g2_decap_8 FILLER_4_120 ();
 sg13g2_decap_8 FILLER_4_127 ();
 sg13g2_decap_8 FILLER_4_134 ();
 sg13g2_decap_8 FILLER_4_141 ();
 sg13g2_decap_8 FILLER_4_148 ();
 sg13g2_decap_8 FILLER_4_155 ();
 sg13g2_decap_4 FILLER_4_162 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_fill_2 FILLER_5_21 ();
 sg13g2_fill_1 FILLER_5_23 ();
 sg13g2_decap_8 FILLER_5_100 ();
 sg13g2_decap_8 FILLER_5_107 ();
 sg13g2_decap_8 FILLER_5_114 ();
 sg13g2_decap_4 FILLER_5_121 ();
 sg13g2_fill_1 FILLER_5_125 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_158 ();
 sg13g2_fill_1 FILLER_5_165 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_10 ();
 sg13g2_decap_8 FILLER_6_17 ();
 sg13g2_fill_2 FILLER_6_24 ();
 sg13g2_fill_1 FILLER_6_26 ();
 sg13g2_fill_2 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_fill_2 FILLER_6_63 ();
 sg13g2_fill_1 FILLER_6_65 ();
 sg13g2_fill_1 FILLER_6_78 ();
 sg13g2_fill_2 FILLER_6_88 ();
 sg13g2_decap_8 FILLER_6_103 ();
 sg13g2_decap_8 FILLER_6_110 ();
 sg13g2_decap_8 FILLER_6_117 ();
 sg13g2_fill_2 FILLER_6_124 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_fill_2 FILLER_6_137 ();
 sg13g2_decap_4 FILLER_6_143 ();
 sg13g2_fill_1 FILLER_6_151 ();
 sg13g2_decap_4 FILLER_6_156 ();
 sg13g2_fill_2 FILLER_6_160 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_4 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_11 ();
 sg13g2_fill_1 FILLER_7_17 ();
 sg13g2_fill_2 FILLER_7_22 ();
 sg13g2_fill_1 FILLER_7_24 ();
 sg13g2_fill_1 FILLER_7_37 ();
 sg13g2_fill_2 FILLER_7_64 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_decap_4 FILLER_7_125 ();
 sg13g2_fill_2 FILLER_7_133 ();
 sg13g2_fill_1 FILLER_7_153 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_15 ();
 sg13g2_decap_4 FILLER_8_34 ();
 sg13g2_fill_2 FILLER_8_47 ();
 sg13g2_fill_2 FILLER_8_57 ();
 sg13g2_fill_1 FILLER_8_64 ();
 sg13g2_fill_1 FILLER_8_83 ();
 sg13g2_decap_8 FILLER_8_92 ();
 sg13g2_decap_8 FILLER_8_99 ();
 sg13g2_fill_1 FILLER_8_106 ();
 sg13g2_fill_2 FILLER_8_115 ();
 sg13g2_fill_1 FILLER_8_142 ();
 sg13g2_decap_4 FILLER_8_160 ();
 sg13g2_fill_2 FILLER_8_164 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_16 ();
 sg13g2_fill_1 FILLER_9_23 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_4 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_99 ();
 sg13g2_fill_2 FILLER_9_106 ();
 sg13g2_fill_2 FILLER_9_121 ();
 sg13g2_fill_2 FILLER_9_136 ();
 sg13g2_fill_1 FILLER_9_143 ();
 sg13g2_decap_4 FILLER_9_151 ();
 sg13g2_fill_2 FILLER_9_163 ();
 sg13g2_fill_1 FILLER_9_165 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_fill_1 FILLER_10_11 ();
 sg13g2_fill_2 FILLER_10_16 ();
 sg13g2_fill_1 FILLER_10_18 ();
 sg13g2_fill_1 FILLER_10_23 ();
 sg13g2_fill_1 FILLER_10_29 ();
 sg13g2_fill_1 FILLER_10_38 ();
 sg13g2_fill_2 FILLER_10_44 ();
 sg13g2_fill_1 FILLER_10_59 ();
 sg13g2_fill_2 FILLER_10_76 ();
 sg13g2_decap_4 FILLER_10_115 ();
 sg13g2_fill_1 FILLER_10_119 ();
 sg13g2_fill_1 FILLER_10_147 ();
 sg13g2_fill_2 FILLER_10_153 ();
 sg13g2_decap_4 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_11 ();
 sg13g2_fill_1 FILLER_11_17 ();
 sg13g2_fill_1 FILLER_11_22 ();
 sg13g2_fill_2 FILLER_11_35 ();
 sg13g2_fill_1 FILLER_11_40 ();
 sg13g2_fill_2 FILLER_11_46 ();
 sg13g2_fill_2 FILLER_11_56 ();
 sg13g2_fill_2 FILLER_11_62 ();
 sg13g2_fill_1 FILLER_11_64 ();
 sg13g2_fill_2 FILLER_11_69 ();
 sg13g2_fill_1 FILLER_11_71 ();
 sg13g2_fill_2 FILLER_11_76 ();
 sg13g2_fill_2 FILLER_11_91 ();
 sg13g2_fill_1 FILLER_11_93 ();
 sg13g2_fill_1 FILLER_11_140 ();
 sg13g2_fill_2 FILLER_11_146 ();
 sg13g2_fill_1 FILLER_11_156 ();
 sg13g2_fill_1 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_fill_1 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_30 ();
 sg13g2_decap_4 FILLER_12_47 ();
 sg13g2_fill_1 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_77 ();
 sg13g2_fill_1 FILLER_12_79 ();
 sg13g2_fill_1 FILLER_12_88 ();
 sg13g2_decap_8 FILLER_12_93 ();
 sg13g2_decap_4 FILLER_12_100 ();
 sg13g2_fill_1 FILLER_12_129 ();
 sg13g2_fill_1 FILLER_12_142 ();
 sg13g2_fill_2 FILLER_12_164 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_30 ();
 sg13g2_fill_2 FILLER_13_40 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_fill_2 FILLER_13_57 ();
 sg13g2_fill_1 FILLER_13_59 ();
 sg13g2_fill_2 FILLER_13_64 ();
 sg13g2_decap_4 FILLER_13_70 ();
 sg13g2_fill_2 FILLER_13_90 ();
 sg13g2_fill_1 FILLER_13_92 ();
 sg13g2_decap_4 FILLER_13_112 ();
 sg13g2_fill_2 FILLER_13_128 ();
 sg13g2_fill_1 FILLER_13_142 ();
 sg13g2_fill_1 FILLER_13_147 ();
 sg13g2_fill_1 FILLER_13_156 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_82 ();
 sg13g2_fill_2 FILLER_14_87 ();
 sg13g2_fill_1 FILLER_14_94 ();
 sg13g2_decap_8 FILLER_14_103 ();
 sg13g2_fill_2 FILLER_14_110 ();
 sg13g2_fill_2 FILLER_14_120 ();
 sg13g2_fill_1 FILLER_14_122 ();
 sg13g2_fill_2 FILLER_14_127 ();
 sg13g2_fill_1 FILLER_14_129 ();
 sg13g2_fill_1 FILLER_14_139 ();
 sg13g2_fill_2 FILLER_14_154 ();
 sg13g2_fill_1 FILLER_14_160 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_4 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_32 ();
 sg13g2_fill_1 FILLER_15_46 ();
 sg13g2_fill_1 FILLER_15_53 ();
 sg13g2_fill_1 FILLER_15_59 ();
 sg13g2_fill_1 FILLER_15_68 ();
 sg13g2_fill_2 FILLER_15_74 ();
 sg13g2_decap_4 FILLER_15_83 ();
 sg13g2_decap_8 FILLER_15_100 ();
 sg13g2_decap_8 FILLER_15_107 ();
 sg13g2_fill_1 FILLER_15_114 ();
 sg13g2_decap_8 FILLER_15_129 ();
 sg13g2_fill_2 FILLER_15_136 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_28 ();
 sg13g2_fill_1 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_51 ();
 sg13g2_fill_1 FILLER_16_62 ();
 sg13g2_fill_1 FILLER_16_86 ();
 sg13g2_decap_8 FILLER_16_95 ();
 sg13g2_decap_4 FILLER_16_102 ();
 sg13g2_fill_1 FILLER_16_106 ();
 sg13g2_decap_8 FILLER_16_111 ();
 sg13g2_decap_4 FILLER_16_118 ();
 sg13g2_fill_2 FILLER_16_122 ();
 sg13g2_fill_2 FILLER_16_138 ();
 sg13g2_fill_1 FILLER_16_152 ();
 sg13g2_fill_1 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_42 ();
 sg13g2_decap_4 FILLER_17_52 ();
 sg13g2_fill_1 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_65 ();
 sg13g2_decap_8 FILLER_17_72 ();
 sg13g2_decap_8 FILLER_17_79 ();
 sg13g2_decap_8 FILLER_17_86 ();
 sg13g2_decap_8 FILLER_17_93 ();
 sg13g2_decap_4 FILLER_17_100 ();
 sg13g2_fill_2 FILLER_17_163 ();
 sg13g2_fill_1 FILLER_17_165 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_fill_2 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_55 ();
 sg13g2_fill_2 FILLER_18_62 ();
 sg13g2_fill_1 FILLER_18_64 ();
 sg13g2_fill_1 FILLER_18_109 ();
 sg13g2_fill_2 FILLER_18_122 ();
 sg13g2_fill_2 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_157 ();
 sg13g2_fill_2 FILLER_18_164 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_4 FILLER_19_46 ();
 sg13g2_fill_1 FILLER_19_102 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_fill_1 FILLER_19_131 ();
 sg13g2_fill_1 FILLER_19_136 ();
 sg13g2_fill_1 FILLER_19_142 ();
 sg13g2_fill_1 FILLER_19_151 ();
 sg13g2_fill_2 FILLER_19_164 ();
endmodule
